BZh91AY&SY4Σ j_�py���������P��r��
 $�e=&��S4��5#@ 4 h jy&T�@ �#   $�PT����40!� ���&L��L �0L�0�D�OF�@�ɔ�z�F��CCOBfS�~�PH�$��H���l6� s�g?���I�I�&�R�J�[cS#a*��1[@H�d�iGic���p���f�AhC.��a�kŽ}�Ls.��ȸ����;#"z9A��0{'R�v���� BS��	%Tk9����߷��� �^�ыM+�sh��J� �&��XH���4����l�kr�,)ޫ�,�^d�	l�óRSX)�i�@���i��,RaJs �LX�t����
�^]3ܡ�!&t��Uo1n��5�ԙiF��54�񲨢�YUE-��7{�@�n��ŕp�ꆆ@��@�����+ܜ�
Ln��W1����/E�@NM�k�&�m^�U�~�~Xo����D�u�ɩ��X'�ő5f�����oL�WL����1�\�3�����B.�hc*��F����HA�x =��dG'>��94{�3�4@��,�x/��aN ��d��m���TO~�B�@|mT5������x?�V�	ёYYJU�5u�jj��,�5%/�"�* #{E�l�J\� j��,d�)´<i w�9�Z�IS�� ℸ���;In���?+��0��fQVk�?I����s��`�h�=Y!y$�3O�f��F	�PBҼ��;�/,GEwЮ��P���(�}��a�Z���������K���N��]Q�!l�B�%�������tA�;�]Ay�i@E� �dGNd �0�B�78�b\PE��8��҅�JXU �3w?�Dm6�3�$�4Y��$CH�8"ԭ[p*�N)���d-�&x�9��Z���P����9�4@i����A�9}���i�
*65x3r�᧶Nd�N�����5��ߊ�Am�of�gt�̇�<-@W$��N5cزQ����o�Y�Yac@i�j��J��U�b4y<t�����0(�ىsf�D�TD�}!O���!w��P���`s&0W`Y���"�(HgQ� 